module tb_top_level;

endmodule
