module video_memory;



endmodule

