`timescale 1ns / 1ps

// Multiplier-Accumulator 
module mac();

endmodule

