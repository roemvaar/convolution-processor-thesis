// Control Unit
//
// Steps:
// 1. At startup, load weights at each processing elements that compose the systolic array
// 2.
//

module control_unit;

endmodule
