// Define n processing elements

module systolic_array;

endmodule

