module tb_mac;

    // Inputs
    reg[] in_a;
    reg[] in_b; 
    
endmodule

