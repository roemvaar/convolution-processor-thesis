`timescale 1ns / 1ps

// Multiplier-Accumulator (MAC)
// The multiply-accumulate operation is a common step that
// computes the product of two numbers and adds that product
// to an accumulator.
// a <- a + (b x c)
module mac();

endmodule

