module proc_elem;

endmodule

