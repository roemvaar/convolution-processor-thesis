// Define n processing elements

module systolic_array (x, k, h);
    input x;
    input k;
    output h;

    parameter DATA_WIDTH = 16;

endmodule
 
