module toplevel;


endmodule

