module tb_systolic_array;

endmodule
