module tb_control_unit;

endmodule
