module tb_video_memory;


endmodule
