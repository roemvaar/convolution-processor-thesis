module systolic_array;
endmodule

