module tb_proc_elem;

endmodule
